version https://git-lfs.github.com/spec/v1
oid sha256:ed773d4d9f2a01b7b866c25cda6961130c65e594f30c1e5b087e1588906f2dac
size 230
